module toSegment(boxRow0,boxRow1,boxRow2,boxRow3,boxColumn,xOuts,yOuts,count);
    input boxRow

endmodule